module clb (
    input [127:0]a , b ,
    output [127:0] c 
);
assign c = a + b ;
    
endmodule